package motion_estimator_test_pkg;
import uvm_pkg::*;
import motion_estimator_env_pkg::*;
import motion_estimator_agent_pkg::*;
 `include "motion_estimator_seq.sv"
 `include "motion_estimator_msb_bits_seq.sv"
 `include "motion_estimator_rf_ffff_sf_ffff_seq.sv"
 `include "motion_estimator_test.sv"
 `include "motion_estimator_rf_msb_bits_test.sv"
 `include "motion_estimator_s1_msb_bits_test.sv"
 `include "motion_estimator_s2_msb_bits_test.sv"
 `include "motion_estimator_rf_ffff_sf_ffff_test.sv"
endpackage
