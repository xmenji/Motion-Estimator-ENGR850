package motion_estimator_env_pkg;
import uvm_pkg::*;
import motion_estimator_agent_pkg::*;
localparam string s_motion_estimator_env_config_id = "tb_top_level_config";
 `include "motion_estimator_virtual_sequencer.sv"
 `include "motion_estimator_env_config.sv"
 `include "motion_estimator_scoreboard.sv"
 `include "motion_estimator_env.sv"
endpackage
