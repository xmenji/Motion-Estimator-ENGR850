//driver, monitor,seq item,sequence are included here . if oyu pas this for
//cmpialtion will take all the required files
package motion_estimator_agent_pkg;
 import uvm_pkg::*;
  `include "motion_estimator_sequence_item.sv"
  `include "motion_estimator_driver.sv"
  `include "motion_estimator_sequencer.sv"
  `include "motion_estimator_cov.sv"
  `include "motion_estimator_monitor.sv"
  `include "motion_estimator_agent.sv"
endpackage 
